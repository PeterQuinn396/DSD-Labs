library verilog;
use verilog.vl_types.all;
entity g07_pop_enable_vlg_vec_tst is
end g07_pop_enable_vlg_vec_tst;
