library verilog;
use verilog.vl_types.all;
entity g07_lab5_testbed_vlg_vec_tst is
end g07_lab5_testbed_vlg_vec_tst;
