library verilog;
use verilog.vl_types.all;
entity g07_debouncer_vlg_check_tst is
    port(
        sig             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g07_debouncer_vlg_check_tst;
