library verilog;
use verilog.vl_types.all;
entity g07_testing_vlg_vec_tst is
end g07_testing_vlg_vec_tst;
