library verilog;
use verilog.vl_types.all;
entity g07_7_segment_decoder_vlg_vec_tst is
end g07_7_segment_decoder_vlg_vec_tst;
