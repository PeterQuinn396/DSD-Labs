library verilog;
use verilog.vl_types.all;
entity g07_computer_FSM_vlg_vec_tst is
end g07_computer_FSM_vlg_vec_tst;
