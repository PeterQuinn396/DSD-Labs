library verilog;
use verilog.vl_types.all;
entity g07_dealer_FSM_vlg_check_tst is
    port(
        stack_enable    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g07_dealer_FSM_vlg_check_tst;
